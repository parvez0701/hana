module test(input d, clk, reset, set, output reg q);
always @(posedge clk or posedge reset or negedge set) 
    if(reset)
	    q <= 0;
	else if(!set)
	    q <= 1;
	else	
        q <= d;
endmodule	
