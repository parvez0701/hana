module test(in, out);
        input wire in;
    output wire out;

// Variable declaration.
    assign  out = in;


endmodule
