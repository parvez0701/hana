module test();

wire synth_net;
wire synth_net_0;
wire synth_net_1;
wire synth_net_2;
wire synth_net_3;
wire synth_net_4;
wire synth_net_5;
wire synth_net_6;
wire synth_net_7;
wire synth_net_8;
wire synth_net_9;
wire synth_net_10;
wire synth_net_11;
wire synth_net_12;
wire synth_net_13;
wire synth_net_14;
wire synth_net_15;
wire synth_net_16;
wire synth_net_17;
wire synth_net_18;
wire synth_net_19;
wire synth_net_20;
wire synth_net_21;
wire synth_net_22;
wire synth_net_23;
wire synth_net_24;
wire synth_net_25;
wire synth_net_26;
wire synth_net_27;
wire synth_net_28;
reg [1:0] A;
reg [1:0] B;
reg [1:0] AB_AND;
reg [1:0] AB_OR;
reg [1:0] AB_XOR;
reg ab_and;
AND_2_1 synth_AND(.OUT(synth_net), .IN({A[1], B[1]}));
AND_2_1 synth_AND_0(.OUT(synth_net_0), .IN({A[0], B[0]}));
BUF_1_1 synth_BUF(.OUT(synth_net_1), .IN(synth_net));
VCC_0_1 synth_VCC(.OUT(synth_net_2));
BUF_1_1 synth_BUF_0(.OUT(synth_net_3), .IN(synth_net_0));
VCC_0_1 synth_VCC_0(.OUT(synth_net_4));
OR_2_1 synth_OR(.OUT(synth_net_5), .IN({A[1], B[1]}));
OR_2_1 synth_OR_0(.OUT(synth_net_6), .IN({A[0], B[0]}));
BUF_1_1 synth_BUF_1(.OUT(synth_net_7), .IN(synth_net_5));
VCC_0_1 synth_VCC_1(.OUT(synth_net_8));
BUF_1_1 synth_BUF_2(.OUT(synth_net_9), .IN(synth_net_6));
VCC_0_1 synth_VCC_2(.OUT(synth_net_10));
XOR_2_1 synth_XOR(.OUT(synth_net_11), .IN({A[1], B[1]}));
XOR_2_1 synth_XOR_0(.OUT(synth_net_12), .IN({A[0], B[0]}));
BUF_1_1 synth_BUF_3(.OUT(synth_net_13), .IN(synth_net_11));
VCC_0_1 synth_VCC_3(.OUT(synth_net_14));
BUF_1_1 synth_BUF_4(.OUT(synth_net_15), .IN(synth_net_12));
VCC_0_1 synth_VCC_4(.OUT(synth_net_16));
AND_2_1 synth_AND_1(.OUT(synth_net_17), .IN({synth_net_13, synth_net_14}));
AND_2_1 synth_AND_2(.OUT(synth_net_18), .IN({synth_net_15, synth_net_16}));
AND_2_1 synth_AND_3(.OUT(synth_net_19), .IN({synth_net_7, synth_net_8}));
AND_2_1 synth_AND_4(.OUT(synth_net_20), .IN({synth_net_9, synth_net_10}));
AND_2_1 synth_AND_5(.OUT(synth_net_21), .IN({synth_net_1, synth_net_2}));
AND_2_1 synth_AND_6(.OUT(synth_net_22), .IN({synth_net_3, synth_net_4}));
AND_2_1 synth_AND_7(.OUT(synth_net_23), .IN({synth_net_21, synth_net_2}));
BUF_1_1 synth_BUF_5(.OUT(AB_AND[1]), .IN(synth_net_23));
AND_2_1 synth_AND_8(.OUT(synth_net_24), .IN({synth_net_22, synth_net_4}));
BUF_1_1 synth_BUF_6(.OUT(AB_AND[0]), .IN(synth_net_24));
AND_2_1 synth_AND_9(.OUT(synth_net_25), .IN({synth_net_19, synth_net_8}));
BUF_1_1 synth_BUF_7(.OUT(AB_OR[1]), .IN(synth_net_25));
AND_2_1 synth_AND_10(.OUT(synth_net_26), .IN({synth_net_20, synth_net_10}));
BUF_1_1 synth_BUF_8(.OUT(AB_OR[0]), .IN(synth_net_26));
AND_2_1 synth_AND_11(.OUT(synth_net_27), .IN({synth_net_17, synth_net_14}));
BUF_1_1 synth_BUF_9(.OUT(AB_XOR[1]), .IN(synth_net_27));
AND_2_1 synth_AND_12(.OUT(synth_net_28), .IN({synth_net_18, synth_net_16}));
BUF_1_1 synth_BUF_10(.OUT(AB_XOR[0]), .IN(synth_net_28));
endmodule
