module test (output [1:0] out);
assign out = 2'sb11;
endmodule
