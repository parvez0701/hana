module test(input in1, in2, in3, in4, in5, in6,  
    in7, in8, in9, in10, in11, in12, output out1, out2);
assign out1 = in1 & in2 & in3 & in4 & in5 & in6;
assign out2 = in7 | in8 | in9 | in10 | in11 | in12;
endmodule
