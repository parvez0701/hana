module test();

reg reg1;
reg [1:0] reg2;
reg [1:0] reg3;
reg [9:0] reg4;
endmodule
