module test();
reg reg1;
reg [1:0] reg2;
reg reg3 [1:0];
reg [1:0] reg4 [0:4];
endmodule
