
module LIBMOD1();
endmodule

module LIBMOD();
LIBMOD1 L1();
endmodule
