module test();
    wire w;
    
// Variable declaration.


endmodule
