module test();
wire wire1;
wire [1:0] wire2;
wire wire3 [1:0];
wire [1:0] wire4 [0:4];
endmodule
