module test();

task check_result (input [63:0] result,
					input [63:0] expected,
					output	OK);

	begin
	end

endtask

function integer fp_alu(input reg r1);

begin
end
endfunction

endmodule
					
