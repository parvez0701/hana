module test(in, out, io);

input wire in;
output wire out;
inout wire io;
endmodule
