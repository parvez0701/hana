module test();
    
// Variable declaration.


    task check_result;
    input  [63:0] result ;
    input  [63:0] expected ;
    output  OK;

// Variable declaration.
    begin
    end
    endtask
    function integer fp_alu;
    input reg r1;

// Variable declaration.
    integer  fp_alu;
    begin
    end
    endfunction

endmodule
