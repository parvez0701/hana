module adder(	output	reg		[31:0]	sum [1:0],
				output	reg				co,
				input	wire	[31:0]	a,
				input	wire	[31:0]	b,
				input	wire			ci);
endmodule	
