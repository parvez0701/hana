module test();
integer integer1;
integer  integer2;
integer integer3 [1:0];
integer integer4 [1:0][0:4];
endmodule
