module test(in1, in2, out);
        input wire in1;
    input wire in2;
    output wire out;

// Variable declaration.
    assign  out = in1;


endmodule
