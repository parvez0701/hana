module test(input in, output out);
wire w;
and(w, w, w);
endmodule
