module test(in, out);

input wire [7:0]in;
output wire [7:0]out;
wire [7:0]byte0;
wire [7:0]byte2;
wire [7:0]byte3;
wire [7:0]byte4;
wire synth_net;
wire synth_net_0;
wire synth_net_1;
wire synth_net_2;
wire synth_net_3;
wire synth_net_4;
wire synth_net_5;
wire synth_net_6;
wire synth_net_7;
wire synth_net_8;
wire synth_net_9;
wire synth_net_10;
wire synth_net_11;
wire synth_net_12;
wire synth_net_13;
wire synth_net_14;
wire synth_net_15;
wire synth_net_16;
wire synth_net_17;
wire synth_net_18;
wire synth_net_19;
wire synth_net_20;
wire synth_net_21;
wire synth_net_22;
wire synth_net_23;
wire synth_net_24;
wire synth_net_25;
wire synth_net_26;
wire synth_net_27;
wire synth_net_28;
wire synth_net_29;
wire synth_net_30;
wire synth_net_31;
wire synth_net_32;
wire synth_net_33;
wire synth_net_34;
wire synth_net_35;
wire synth_net_36;
wire synth_net_37;
wire synth_net_38;
reg [255:0] data1;
reg [0:255] data2;
reg [7:0] byte1;
reg signed [31:0] i;
BUF_1_1 synth_BUF(.OUT(out[5]), .IN(in[3]));
BUF_1_1 synth_BUF_0(.OUT(out[4]), .IN(in[2]));
BUF_1_1 synth_BUF_1(.OUT(out[3]), .IN(in[1]));
BUF_1_1 synth_BUF_2(.OUT(out[2]), .IN(in[0]));
BUF_1_1 synth_BUF_3(.OUT(byte0[7]), .IN(data1[30]));
BUF_1_1 synth_BUF_4(.OUT(byte0[6]), .IN(data1[29]));
BUF_1_1 synth_BUF_5(.OUT(byte0[5]), .IN(data1[28]));
BUF_1_1 synth_BUF_6(.OUT(byte0[4]), .IN(data1[27]));
BUF_1_1 synth_BUF_7(.OUT(byte0[3]), .IN(data1[26]));
BUF_1_1 synth_BUF_8(.OUT(byte0[2]), .IN(data1[25]));
BUF_1_1 synth_BUF_9(.OUT(byte0[1]), .IN(data1[24]));
BUF_1_1 synth_BUF_10(.OUT(byte0[0]), .IN(data1[23]));
BUF_1_1 synth_BUF_11(.OUT(byte2[7]), .IN(data1[31]));
BUF_1_1 synth_BUF_12(.OUT(byte2[6]), .IN(data1[30]));
BUF_1_1 synth_BUF_13(.OUT(byte2[5]), .IN(data1[29]));
BUF_1_1 synth_BUF_14(.OUT(byte2[4]), .IN(data1[28]));
BUF_1_1 synth_BUF_15(.OUT(byte2[3]), .IN(data1[27]));
BUF_1_1 synth_BUF_16(.OUT(byte2[2]), .IN(data1[26]));
BUF_1_1 synth_BUF_17(.OUT(byte2[1]), .IN(data1[25]));
BUF_1_1 synth_BUF_18(.OUT(byte2[0]), .IN(data1[24]));
BUF_1_1 synth_BUF_19(.OUT(byte3[7]), .IN(data2[24]));
BUF_1_1 synth_BUF_20(.OUT(byte3[6]), .IN(data2[25]));
BUF_1_1 synth_BUF_21(.OUT(byte3[5]), .IN(data2[26]));
BUF_1_1 synth_BUF_22(.OUT(byte3[4]), .IN(data2[27]));
BUF_1_1 synth_BUF_23(.OUT(byte3[3]), .IN(data2[28]));
BUF_1_1 synth_BUF_24(.OUT(byte3[2]), .IN(data2[29]));
BUF_1_1 synth_BUF_25(.OUT(byte3[1]), .IN(data2[30]));
BUF_1_1 synth_BUF_26(.OUT(byte3[0]), .IN(data2[31]));
BUF_1_1 synth_BUF_27(.OUT(byte4[7]), .IN(data2[25]));
BUF_1_1 synth_BUF_28(.OUT(byte4[6]), .IN(data2[26]));
BUF_1_1 synth_BUF_29(.OUT(byte4[5]), .IN(data2[27]));
BUF_1_1 synth_BUF_30(.OUT(byte4[4]), .IN(data2[28]));
BUF_1_1 synth_BUF_31(.OUT(byte4[3]), .IN(data2[29]));
BUF_1_1 synth_BUF_32(.OUT(byte4[2]), .IN(data2[30]));
BUF_1_1 synth_BUF_33(.OUT(byte4[1]), .IN(data2[31]));
BUF_1_1 synth_BUF_34(.OUT(byte4[0]), .IN(data2[32]));
BUF_1_1 synth_BUF_35(.OUT(synth_net), .IN(data1[7]));
VCC_0_1 synth_VCC(.OUT(synth_net_0));
BUF_1_1 synth_BUF_36(.OUT(synth_net_1), .IN(data1[6]));
VCC_0_1 synth_VCC_0(.OUT(synth_net_2));
BUF_1_1 synth_BUF_37(.OUT(synth_net_3), .IN(data1[5]));
VCC_0_1 synth_VCC_1(.OUT(synth_net_4));
BUF_1_1 synth_BUF_38(.OUT(synth_net_5), .IN(data1[4]));
VCC_0_1 synth_VCC_2(.OUT(synth_net_6));
BUF_1_1 synth_BUF_39(.OUT(synth_net_7), .IN(data1[3]));
VCC_0_1 synth_VCC_3(.OUT(synth_net_8));
BUF_1_1 synth_BUF_40(.OUT(synth_net_9), .IN(data1[2]));
VCC_0_1 synth_VCC_4(.OUT(synth_net_10));
BUF_1_1 synth_BUF_41(.OUT(synth_net_11), .IN(data1[1]));
VCC_0_1 synth_VCC_5(.OUT(synth_net_12));
BUF_1_1 synth_BUF_42(.OUT(synth_net_13), .IN(data1[0]));
VCC_0_1 synth_VCC_6(.OUT(synth_net_14));
BUF_1_1 synth_BUF_43(.OUT(synth_net_15), .IN(data1[15]));
VCC_0_1 synth_VCC_7(.OUT(synth_net_16));
BUF_1_1 synth_BUF_44(.OUT(synth_net_17), .IN(data1[14]));
VCC_0_1 synth_VCC_8(.OUT(synth_net_18));
BUF_1_1 synth_BUF_45(.OUT(synth_net_19), .IN(data1[13]));
VCC_0_1 synth_VCC_9(.OUT(synth_net_20));
BUF_1_1 synth_BUF_46(.OUT(synth_net_21), .IN(data1[12]));
VCC_0_1 synth_VCC_10(.OUT(synth_net_22));
BUF_1_1 synth_BUF_47(.OUT(synth_net_23), .IN(data1[11]));
VCC_0_1 synth_VCC_11(.OUT(synth_net_24));
BUF_1_1 synth_BUF_48(.OUT(synth_net_25), .IN(data1[10]));
VCC_0_1 synth_VCC_12(.OUT(synth_net_26));
BUF_1_1 synth_BUF_49(.OUT(synth_net_27), .IN(data1[9]));
VCC_0_1 synth_VCC_13(.OUT(synth_net_28));
BUF_1_1 synth_BUF_50(.OUT(synth_net_29), .IN(data1[8]));
VCC_0_1 synth_VCC_14(.OUT(synth_net_30));
AND_2_1 synth_AND(.OUT(synth_net_31), .IN({synth_net_15, synth_net_16}));
BUF_1_1 synth_BUF_51(.OUT(byte1[7]), .IN(synth_net_31));
AND_2_1 synth_AND_0(.OUT(synth_net_32), .IN({synth_net_17, synth_net_18}));
BUF_1_1 synth_BUF_52(.OUT(byte1[6]), .IN(synth_net_32));
AND_2_1 synth_AND_1(.OUT(synth_net_33), .IN({synth_net_19, synth_net_20}));
BUF_1_1 synth_BUF_53(.OUT(byte1[5]), .IN(synth_net_33));
AND_2_1 synth_AND_2(.OUT(synth_net_34), .IN({synth_net_21, synth_net_22}));
BUF_1_1 synth_BUF_54(.OUT(byte1[4]), .IN(synth_net_34));
AND_2_1 synth_AND_3(.OUT(synth_net_35), .IN({synth_net_23, synth_net_24}));
BUF_1_1 synth_BUF_55(.OUT(byte1[3]), .IN(synth_net_35));
AND_2_1 synth_AND_4(.OUT(synth_net_36), .IN({synth_net_25, synth_net_26}));
BUF_1_1 synth_BUF_56(.OUT(byte1[2]), .IN(synth_net_36));
AND_2_1 synth_AND_5(.OUT(synth_net_37), .IN({synth_net_27, synth_net_28}));
BUF_1_1 synth_BUF_57(.OUT(byte1[1]), .IN(synth_net_37));
AND_2_1 synth_AND_6(.OUT(synth_net_38), .IN({synth_net_29, synth_net_30}));
BUF_1_1 synth_BUF_58(.OUT(byte1[0]), .IN(synth_net_38));
endmodule
