module test(out2, io1, io2, in2, out1, in1);

output wire [0:1]out2;
inout wire [1:0]io1;
inout wire [0:1]io2;
input wire [0:1]in2;
output wire [1:0]out1;
input wire [1:0]in1;
endmodule
