module ahmad();
    // Parameter declarations.
    parameter signed [31:0]param = 10;
wire w;
    
// Variable declaration.
    assign  w = 10;


endmodule
