module test(in, out);

input wire in;
output wire out;
assign out = 0;
endmodule
