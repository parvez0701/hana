module test();
    
// Variable declaration.


endmodule
