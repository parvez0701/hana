module test(output out, input in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21);
assign out = in1 ~^ in2 ~^ in3 ~^ in4 ~^ in5 ~^ in6 ~^ in7 ~^ in8 ~^ in9 ~^ in10 ~^ in11 ~^ in12 ~^ in13 ~^ in14 ~^ in15 ~^ in16 ~^ in17 ~^ in18 ~^ in19 ~^ in20 ~^ in21;
endmodule
