module test(input IN, SHIFT, output OUT);

assign OUT = IN << SHIFT;
endmodule
