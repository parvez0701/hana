module test();
integer integer1;
integer  integer2;
integer integer3 [1:0];
integer integer4 [1:0][0:4];
endmodule

module test1();
real integer1;
real  integer2;
real integer3 [1:0];
real integer4 [1:0][0:4];
endmodule
