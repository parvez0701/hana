
module test ()
endmodule
