module test(out);
        output wire [1:0] out ;

// Variable declaration.
    assign  out = 2'sb11;


endmodule
