module adder (a, b, sum);
	input signed [63:0] a, b;
	output signed sum;
	wire [63:0] a, b;
	reg [63:0] sum;
endmodule
