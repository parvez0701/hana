module test(output out, input in1, in2, in3, in4);

nand mynand(out,  in1, in2, in3, in4 );

endmodule
