module FlipFlop(clk, cs, ns);

input wire clk;
input wire [31:0]cs;
output wire [31:0]ns;
wire synth_net_0;
wire synth_net_2;
wire synth_net_4;
wire synth_net_6;
wire synth_net_8;
wire synth_net_10;
wire synth_net_12;
wire synth_net_14;
wire synth_net_16;
wire synth_net_18;
wire synth_net_20;
wire synth_net_22;
wire synth_net_24;
wire synth_net_26;
wire synth_net_28;
wire synth_net_30;
wire synth_net_32;
wire synth_net_34;
wire synth_net_36;
wire synth_net_38;
wire synth_net_40;
wire synth_net_42;
wire synth_net_44;
wire synth_net_46;
wire synth_net_48;
wire synth_net_50;
wire synth_net_52;
wire synth_net_54;
wire synth_net_56;
wire synth_net_58;
wire synth_net_60;
wire synth_net_62;
wire synth_net_63;
wire synth_net_64;
wire synth_net_65;
wire synth_net_66;
wire synth_net_67;
wire synth_net_68;
wire synth_net_69;
wire synth_net_70;
wire synth_net_71;
wire synth_net_72;
wire synth_net_73;
wire synth_net_74;
wire synth_net_75;
wire synth_net_76;
wire synth_net_77;
wire synth_net_78;
wire synth_net_79;
wire synth_net_80;
wire synth_net_81;
wire synth_net_82;
wire synth_net_83;
wire synth_net_84;
wire synth_net_85;
wire synth_net_86;
wire synth_net_87;
wire synth_net_88;
wire synth_net_89;
wire synth_net_90;
wire synth_net_91;
wire synth_net_92;
wire synth_net_93;
wire synth_net_94;
reg signed [31:0] is;
VCC_0_1 synth_VCC(.OUT(synth_net_0));
VCC_0_1 synth_VCC_0(.OUT(synth_net_2));
VCC_0_1 synth_VCC_1(.OUT(synth_net_4));
VCC_0_1 synth_VCC_2(.OUT(synth_net_6));
VCC_0_1 synth_VCC_3(.OUT(synth_net_8));
VCC_0_1 synth_VCC_4(.OUT(synth_net_10));
VCC_0_1 synth_VCC_5(.OUT(synth_net_12));
VCC_0_1 synth_VCC_6(.OUT(synth_net_14));
VCC_0_1 synth_VCC_7(.OUT(synth_net_16));
VCC_0_1 synth_VCC_8(.OUT(synth_net_18));
VCC_0_1 synth_VCC_9(.OUT(synth_net_20));
VCC_0_1 synth_VCC_10(.OUT(synth_net_22));
VCC_0_1 synth_VCC_11(.OUT(synth_net_24));
VCC_0_1 synth_VCC_12(.OUT(synth_net_26));
VCC_0_1 synth_VCC_13(.OUT(synth_net_28));
VCC_0_1 synth_VCC_14(.OUT(synth_net_30));
VCC_0_1 synth_VCC_15(.OUT(synth_net_32));
VCC_0_1 synth_VCC_16(.OUT(synth_net_34));
VCC_0_1 synth_VCC_17(.OUT(synth_net_36));
VCC_0_1 synth_VCC_18(.OUT(synth_net_38));
VCC_0_1 synth_VCC_19(.OUT(synth_net_40));
VCC_0_1 synth_VCC_20(.OUT(synth_net_42));
VCC_0_1 synth_VCC_21(.OUT(synth_net_44));
VCC_0_1 synth_VCC_22(.OUT(synth_net_46));
VCC_0_1 synth_VCC_23(.OUT(synth_net_48));
VCC_0_1 synth_VCC_24(.OUT(synth_net_50));
VCC_0_1 synth_VCC_25(.OUT(synth_net_52));
VCC_0_1 synth_VCC_26(.OUT(synth_net_54));
VCC_0_1 synth_VCC_27(.OUT(synth_net_56));
VCC_0_1 synth_VCC_28(.OUT(synth_net_58));
VCC_0_1 synth_VCC_29(.OUT(synth_net_60));
VCC_0_1 synth_VCC_30(.OUT(synth_net_62));
AND_2_1 synth_AND(.OUT(synth_net_63), .IN({synth_net, synth_net_0}));
FF_2_1 synth_FF(.Q(ns[31]), .D(synth_net_63), .CLK(clk));
AND_2_1 synth_AND_0(.OUT(synth_net_64), .IN({synth_net_1, synth_net_2}));
FF_2_1 synth_FF_0(.Q(ns[30]), .D(synth_net_64), .CLK(clk));
AND_2_1 synth_AND_1(.OUT(synth_net_65), .IN({synth_net_3, synth_net_4}));
FF_2_1 synth_FF_1(.Q(ns[29]), .D(synth_net_65), .CLK(clk));
AND_2_1 synth_AND_2(.OUT(synth_net_66), .IN({synth_net_5, synth_net_6}));
FF_2_1 synth_FF_2(.Q(ns[28]), .D(synth_net_66), .CLK(clk));
AND_2_1 synth_AND_3(.OUT(synth_net_67), .IN({synth_net_7, synth_net_8}));
FF_2_1 synth_FF_3(.Q(ns[27]), .D(synth_net_67), .CLK(clk));
AND_2_1 synth_AND_4(.OUT(synth_net_68), .IN({synth_net_9, synth_net_10}));
FF_2_1 synth_FF_4(.Q(ns[26]), .D(synth_net_68), .CLK(clk));
AND_2_1 synth_AND_5(.OUT(synth_net_69), .IN({synth_net_11, synth_net_12}));
FF_2_1 synth_FF_5(.Q(ns[25]), .D(synth_net_69), .CLK(clk));
AND_2_1 synth_AND_6(.OUT(synth_net_70), .IN({synth_net_13, synth_net_14}));
FF_2_1 synth_FF_6(.Q(ns[24]), .D(synth_net_70), .CLK(clk));
AND_2_1 synth_AND_7(.OUT(synth_net_71), .IN({synth_net_15, synth_net_16}));
FF_2_1 synth_FF_7(.Q(ns[23]), .D(synth_net_71), .CLK(clk));
AND_2_1 synth_AND_8(.OUT(synth_net_72), .IN({synth_net_17, synth_net_18}));
FF_2_1 synth_FF_8(.Q(ns[22]), .D(synth_net_72), .CLK(clk));
AND_2_1 synth_AND_9(.OUT(synth_net_73), .IN({synth_net_19, synth_net_20}));
FF_2_1 synth_FF_9(.Q(ns[21]), .D(synth_net_73), .CLK(clk));
AND_2_1 synth_AND_10(.OUT(synth_net_74), .IN({synth_net_21, synth_net_22}));
FF_2_1 synth_FF_10(.Q(ns[20]), .D(synth_net_74), .CLK(clk));
AND_2_1 synth_AND_11(.OUT(synth_net_75), .IN({synth_net_23, synth_net_24}));
FF_2_1 synth_FF_11(.Q(ns[19]), .D(synth_net_75), .CLK(clk));
AND_2_1 synth_AND_12(.OUT(synth_net_76), .IN({synth_net_25, synth_net_26}));
FF_2_1 synth_FF_12(.Q(ns[18]), .D(synth_net_76), .CLK(clk));
AND_2_1 synth_AND_13(.OUT(synth_net_77), .IN({synth_net_27, synth_net_28}));
FF_2_1 synth_FF_13(.Q(ns[17]), .D(synth_net_77), .CLK(clk));
AND_2_1 synth_AND_14(.OUT(synth_net_78), .IN({synth_net_29, synth_net_30}));
FF_2_1 synth_FF_14(.Q(ns[16]), .D(synth_net_78), .CLK(clk));
AND_2_1 synth_AND_15(.OUT(synth_net_79), .IN({synth_net_31, synth_net_32}));
FF_2_1 synth_FF_15(.Q(ns[15]), .D(synth_net_79), .CLK(clk));
AND_2_1 synth_AND_16(.OUT(synth_net_80), .IN({synth_net_33, synth_net_34}));
FF_2_1 synth_FF_16(.Q(ns[14]), .D(synth_net_80), .CLK(clk));
AND_2_1 synth_AND_17(.OUT(synth_net_81), .IN({synth_net_35, synth_net_36}));
FF_2_1 synth_FF_17(.Q(ns[13]), .D(synth_net_81), .CLK(clk));
AND_2_1 synth_AND_18(.OUT(synth_net_82), .IN({synth_net_37, synth_net_38}));
FF_2_1 synth_FF_18(.Q(ns[12]), .D(synth_net_82), .CLK(clk));
AND_2_1 synth_AND_19(.OUT(synth_net_83), .IN({synth_net_39, synth_net_40}));
FF_2_1 synth_FF_19(.Q(ns[11]), .D(synth_net_83), .CLK(clk));
AND_2_1 synth_AND_20(.OUT(synth_net_84), .IN({synth_net_41, synth_net_42}));
FF_2_1 synth_FF_20(.Q(ns[10]), .D(synth_net_84), .CLK(clk));
AND_2_1 synth_AND_21(.OUT(synth_net_85), .IN({synth_net_43, synth_net_44}));
FF_2_1 synth_FF_21(.Q(ns[9]), .D(synth_net_85), .CLK(clk));
AND_2_1 synth_AND_22(.OUT(synth_net_86), .IN({synth_net_45, synth_net_46}));
FF_2_1 synth_FF_22(.Q(ns[8]), .D(synth_net_86), .CLK(clk));
AND_2_1 synth_AND_23(.OUT(synth_net_87), .IN({synth_net_47, synth_net_48}));
FF_2_1 synth_FF_23(.Q(ns[7]), .D(synth_net_87), .CLK(clk));
AND_2_1 synth_AND_24(.OUT(synth_net_88), .IN({synth_net_49, synth_net_50}));
FF_2_1 synth_FF_24(.Q(ns[6]), .D(synth_net_88), .CLK(clk));
AND_2_1 synth_AND_25(.OUT(synth_net_89), .IN({synth_net_51, synth_net_52}));
FF_2_1 synth_FF_25(.Q(ns[5]), .D(synth_net_89), .CLK(clk));
AND_2_1 synth_AND_26(.OUT(synth_net_90), .IN({synth_net_53, synth_net_54}));
FF_2_1 synth_FF_26(.Q(ns[4]), .D(synth_net_90), .CLK(clk));
AND_2_1 synth_AND_27(.OUT(synth_net_91), .IN({synth_net_55, synth_net_56}));
FF_2_1 synth_FF_27(.Q(ns[3]), .D(synth_net_91), .CLK(clk));
AND_2_1 synth_AND_28(.OUT(synth_net_92), .IN({synth_net_57, synth_net_58}));
FF_2_1 synth_FF_28(.Q(ns[2]), .D(synth_net_92), .CLK(clk));
AND_2_1 synth_AND_29(.OUT(synth_net_93), .IN({synth_net_59, synth_net_60}));
FF_2_1 synth_FF_29(.Q(ns[1]), .D(synth_net_93), .CLK(clk));
AND_2_1 synth_AND_30(.OUT(synth_net_94), .IN({synth_net_61, synth_net_62}));
FF_2_1 synth_FF_30(.Q(ns[0]), .D(synth_net_94), .CLK(clk));
endmodule
