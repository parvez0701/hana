module test(in, out, io);
`include in.v
`include out.v

`include assign1.v

endmodule
