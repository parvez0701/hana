module test(a, b, c, d, z);

input wire a;
input wire b;
input wire c;
input wire d;
output reg z;
wire synth_net_0;
wire synth_net_1;
wire synth_net_3;
wire synth_net_5;
wire synth_net_6;
wire synth_net_8;
wire synth_net_9;
wire synth_net_11;
wire synth_net_13;
wire synth_net_14;
wire synth_net_15;
wire synth_net_16;
reg temp1;
reg temp2;
reg synth_reg;
reg synth_reg_0;
XOR_2_1 synth_XOR(.OUT(synth_net_0), .IN({a, b}));
VCC_0_1 synth_VCC(.OUT(synth_net_1));
VCC_0_1 synth_VCC_0(.OUT(synth_net_3));
XOR_2_1 synth_XOR_0(.OUT(synth_net_5), .IN({c, d}));
VCC_0_1 synth_VCC_1(.OUT(synth_net_6));
VCC_0_1 synth_VCC_2(.OUT(synth_net_8));
XOR_2_1 synth_XOR_1(.OUT(synth_net_9), .IN({synth_reg, synth_reg_0}));
VCC_0_1 synth_VCC_3(.OUT(synth_net_11));
AND_2_1 synth_AND(.OUT(z), .IN({synth_net_10, synth_net_11}));
AND_2_1 synth_AND_0(.OUT(synth_net_13), .IN({synth_net_7, synth_net_8}));
AND_2_1 synth_AND_1(.OUT(synth_net_14), .IN({synth_net_5, synth_net_6}));
BUF_1_1 synth_BUF_6(.OUT(temp2), .IN(synth_net_14));
AND_2_1 synth_AND_2(.OUT(synth_net_15), .IN({synth_net_2, synth_net_3}));
AND_2_1 synth_AND_3(.OUT(synth_net_16), .IN({synth_net_0, synth_net_1}));
BUF_1_1 synth_BUF_8(.OUT(temp1), .IN(synth_net_16));
endmodule
