module test(in, out, io);
        input wire in;
    output wire out;
    inout wire io;

// Variable declaration.
    assign  out = in;
    assign  io = in;


endmodule
