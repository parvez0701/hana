module test(out, in);

output wire out;
input wire in;
assign out = (+in);
endmodule
