module adder(sum, co, a, b, ci);
    // Parameter declarations.
    parameter signed [31:0]MSB = 32;
    parameter signed [31:0]LSB = 0;
    output reg [MSB:LSB] sum ;
    output reg co;
    input wire [MSB:LSB] a ;
    input wire [MSB:LSB] b ;
    input wire ci;

// Variable declaration.


endmodule
