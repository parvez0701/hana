module test(in, out);

input wire in;
output wire out;
assign out = (in+in);
assign out = 0;
endmodule
