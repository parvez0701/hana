module test(in, out, io, vin, vout, vio);
        input wire in;
    output wire out;
    inout wire io;
    input wire [3:0] vin ;
    output wire [3:0] vout ;
    inout wire [0:3] vio ;

// Variable declaration.


endmodule
