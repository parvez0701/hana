module test();
reg myreg;
integer myvar;
task check_result (input [63:0] result,
					input [63:0] expected,
					output	OK);
					reg myreg;

	begin
	end

endtask

function integer fp_alu(input reg r1);
reg myvar;
begin
	myvar = myvar + 1;
end
endfunction

endmodule
					
