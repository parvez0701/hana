module ADD1(sum, co, a, b, ci);
	output 	reg	[31:0]	sum = 0;
	output	reg			co = 0;
	input wire [31:0]	a, b;
	input wire ci;
endmodule
