
module LIBMOD();
endmodule
