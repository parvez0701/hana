module adder(a, b, sum);
        input wire signed [63:0] a ;
    input wire signed [63:0] b ;
    output reg signed [63:0] sum ;

// Variable declaration.


endmodule
