`define X 4
module test(input in, output out);

`ifdef Y               
assign out = in;
`endif

endmodule

